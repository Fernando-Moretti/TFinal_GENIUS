module MUX4X1_1bit (
    input [1:0] sel,        // Sinal de seleção de 2 bits (00, 01, 10, 11)
    input in0,             // Entrada 0 (1 bit)
    input in1,             // Entrada 1 (1 bit)
    input in2,             // Entrada 2 (1 bit)
    input in3,             // Entrada 3 (1 bit)
    output reg out        // Saída (1 bit)
);

    always @(*) begin
        case (sel)
            2'b00: out = in0;
            2'b01: out = in1;
            2'b10: out = in2;
            2'b11: out = in3;
            default: out = 1'b0;  // Valor 'x' para caso default (opcional)
        endcase
    end

endmodule